// Comments and desciption of modules have been deliberately ommitted.
// It is up to the student to document and describe the system.

module IF_PC_Add(
		    input [31:0]  PC_IF,
		    output [31:0] PC_Plus_4_IF
		    );

   assign PC_Plus_4_IF=PC_IF+32'd4;

endmodule // IF_PC_Add




   
   
