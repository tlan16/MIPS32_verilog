// add the shifted address offset and PC_Plus_4 from ID stage

module ID_PC_Add(
		 input [31:0]  PC_Plus_4_ID, // actually from ID stage
		 input [31:0]  Instruction_Shift_Left_2_ID,
		 output [31:0] Branch_Dest_ID
		 );

   assign Branch_Dest_ID = PC_Plus_4_ID + Instruction_Shift_Left_2_ID;

endmodule // EX_PC_Add





   
   
