library verilog;
use verilog.vl_types.all;
entity \testbench.v\ is
end \testbench.v\;
