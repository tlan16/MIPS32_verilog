library verilog;
use verilog.vl_types.all;
entity MIPS32_vlg_vec_tst is
end MIPS32_vlg_vec_tst;
