// Comments and desciption of modules have been deliberately ommitted.
// It is up to the student to document and describe the system.

module MEM_Branch_AND(
		      input Branch_MEM,
		      input  Zero_MEM,
		      output PCSrc_MEM
		      );

   assign PCSrc_MEM = Branch_MEM & Zero_MEM;

endmodule // MEM_Branch_AND




   
   
